../vhdl/seven_segment.vhd