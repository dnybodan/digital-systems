../uart_receiver/tx.sv