../uart_receiver/debounce.sv